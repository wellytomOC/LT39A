module Entrada (
    input wire clock
);
    
endmodule