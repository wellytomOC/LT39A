module Sistema (
    input wire clock50MHz, clock1Hz, reset,

    input wire dav,
    input wire[3:0] KeypadData,

    input wire[3:0] AddressIn,
    input wire RWin,

    output wire[3:0] DataOut

);


    
endmodule